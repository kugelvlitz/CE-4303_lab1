
module cpuqsys (
	clk_clk,
	reset_reset_n,
	pio_continue_0_external_connection_export,
	pio_leds_0_external_connection_export);	

	input		clk_clk;
	input		reset_reset_n;
	input		pio_continue_0_external_connection_export;
	output	[7:0]	pio_leds_0_external_connection_export;
endmodule
