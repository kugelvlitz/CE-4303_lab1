// cpuqsys.v

// Generated using ACDS version 20.1 711

`timescale 1 ps / 1 ps
module cpuqsys (
		input  wire        clk_clk,                                     //                                  clk.clk
		output wire [13:0] new_sdram_controller_0_wire_addr,            //          new_sdram_controller_0_wire.addr
		output wire [1:0]  new_sdram_controller_0_wire_ba,              //                                     .ba
		output wire        new_sdram_controller_0_wire_cas_n,           //                                     .cas_n
		output wire        new_sdram_controller_0_wire_cke,             //                                     .cke
		output wire        new_sdram_controller_0_wire_cs_n,            //                                     .cs_n
		inout  wire [31:0] new_sdram_controller_0_wire_dq,              //                                     .dq
		output wire [3:0]  new_sdram_controller_0_wire_dqm,             //                                     .dqm
		output wire        new_sdram_controller_0_wire_ras_n,           //                                     .ras_n
		output wire        new_sdram_controller_0_wire_we_n,            //                                     .we_n
		input  wire        pio_continue_0_external_connection_export,   //   pio_continue_0_external_connection.export
		output wire [6:0]  pio_display1_0_external_connection_export,   //   pio_display1_0_external_connection.export
		output wire [6:0]  pio_display2_0_external_connection_export,   //   pio_display2_0_external_connection.export
		output wire [6:0]  pio_display3_0_external_connection_export,   //   pio_display3_0_external_connection.export
		output wire [6:0]  pio_display4_0_external_connection_export,   //   pio_display4_0_external_connection.export
		output wire [6:0]  pio_display5_0_external_connection_export,   //   pio_display5_0_external_connection.export
		output wire [6:0]  pio_display6_0_external_connection_export,   //   pio_display6_0_external_connection.export
		output wire [7:0]  pio_leds_0_external_connection_export,       //       pio_leds_0_external_connection.export
		input  wire [1:0]  pio_left_right_0_external_connection_export, // pio_left_right_0_external_connection.export
		input  wire [1:0]  pio_up_down_0_external_connection_export,    //    pio_up_down_0_external_connection.export
		input  wire        reset_reset_n                                //                                reset.reset_n
	);

	wire  [31:0] nios2_gen2_0_data_master_readdata;                          // mm_interconnect_0:nios2_gen2_0_data_master_readdata -> nios2_gen2_0:d_readdata
	wire         nios2_gen2_0_data_master_waitrequest;                       // mm_interconnect_0:nios2_gen2_0_data_master_waitrequest -> nios2_gen2_0:d_waitrequest
	wire         nios2_gen2_0_data_master_debugaccess;                       // nios2_gen2_0:debug_mem_slave_debugaccess_to_roms -> mm_interconnect_0:nios2_gen2_0_data_master_debugaccess
	wire  [26:0] nios2_gen2_0_data_master_address;                           // nios2_gen2_0:d_address -> mm_interconnect_0:nios2_gen2_0_data_master_address
	wire   [3:0] nios2_gen2_0_data_master_byteenable;                        // nios2_gen2_0:d_byteenable -> mm_interconnect_0:nios2_gen2_0_data_master_byteenable
	wire         nios2_gen2_0_data_master_read;                              // nios2_gen2_0:d_read -> mm_interconnect_0:nios2_gen2_0_data_master_read
	wire         nios2_gen2_0_data_master_write;                             // nios2_gen2_0:d_write -> mm_interconnect_0:nios2_gen2_0_data_master_write
	wire  [31:0] nios2_gen2_0_data_master_writedata;                         // nios2_gen2_0:d_writedata -> mm_interconnect_0:nios2_gen2_0_data_master_writedata
	wire  [31:0] nios2_gen2_0_instruction_master_readdata;                   // mm_interconnect_0:nios2_gen2_0_instruction_master_readdata -> nios2_gen2_0:i_readdata
	wire         nios2_gen2_0_instruction_master_waitrequest;                // mm_interconnect_0:nios2_gen2_0_instruction_master_waitrequest -> nios2_gen2_0:i_waitrequest
	wire  [26:0] nios2_gen2_0_instruction_master_address;                    // nios2_gen2_0:i_address -> mm_interconnect_0:nios2_gen2_0_instruction_master_address
	wire         nios2_gen2_0_instruction_master_read;                       // nios2_gen2_0:i_read -> mm_interconnect_0:nios2_gen2_0_instruction_master_read
	wire  [31:0] mm_interconnect_0_nios2_gen2_0_debug_mem_slave_readdata;    // nios2_gen2_0:debug_mem_slave_readdata -> mm_interconnect_0:nios2_gen2_0_debug_mem_slave_readdata
	wire         mm_interconnect_0_nios2_gen2_0_debug_mem_slave_waitrequest; // nios2_gen2_0:debug_mem_slave_waitrequest -> mm_interconnect_0:nios2_gen2_0_debug_mem_slave_waitrequest
	wire         mm_interconnect_0_nios2_gen2_0_debug_mem_slave_debugaccess; // mm_interconnect_0:nios2_gen2_0_debug_mem_slave_debugaccess -> nios2_gen2_0:debug_mem_slave_debugaccess
	wire   [8:0] mm_interconnect_0_nios2_gen2_0_debug_mem_slave_address;     // mm_interconnect_0:nios2_gen2_0_debug_mem_slave_address -> nios2_gen2_0:debug_mem_slave_address
	wire         mm_interconnect_0_nios2_gen2_0_debug_mem_slave_read;        // mm_interconnect_0:nios2_gen2_0_debug_mem_slave_read -> nios2_gen2_0:debug_mem_slave_read
	wire   [3:0] mm_interconnect_0_nios2_gen2_0_debug_mem_slave_byteenable;  // mm_interconnect_0:nios2_gen2_0_debug_mem_slave_byteenable -> nios2_gen2_0:debug_mem_slave_byteenable
	wire         mm_interconnect_0_nios2_gen2_0_debug_mem_slave_write;       // mm_interconnect_0:nios2_gen2_0_debug_mem_slave_write -> nios2_gen2_0:debug_mem_slave_write
	wire  [31:0] mm_interconnect_0_nios2_gen2_0_debug_mem_slave_writedata;   // mm_interconnect_0:nios2_gen2_0_debug_mem_slave_writedata -> nios2_gen2_0:debug_mem_slave_writedata
	wire         mm_interconnect_0_timer_0_s1_chipselect;                    // mm_interconnect_0:timer_0_s1_chipselect -> timer_0:chipselect
	wire  [15:0] mm_interconnect_0_timer_0_s1_readdata;                      // timer_0:readdata -> mm_interconnect_0:timer_0_s1_readdata
	wire   [2:0] mm_interconnect_0_timer_0_s1_address;                       // mm_interconnect_0:timer_0_s1_address -> timer_0:address
	wire         mm_interconnect_0_timer_0_s1_write;                         // mm_interconnect_0:timer_0_s1_write -> timer_0:write_n
	wire  [15:0] mm_interconnect_0_timer_0_s1_writedata;                     // mm_interconnect_0:timer_0_s1_writedata -> timer_0:writedata
	wire         mm_interconnect_0_ram_0_s1_chipselect;                      // mm_interconnect_0:ram_0_s1_chipselect -> ram_0:chipselect
	wire  [31:0] mm_interconnect_0_ram_0_s1_readdata;                        // ram_0:readdata -> mm_interconnect_0:ram_0_s1_readdata
	wire  [10:0] mm_interconnect_0_ram_0_s1_address;                         // mm_interconnect_0:ram_0_s1_address -> ram_0:address
	wire   [3:0] mm_interconnect_0_ram_0_s1_byteenable;                      // mm_interconnect_0:ram_0_s1_byteenable -> ram_0:byteenable
	wire         mm_interconnect_0_ram_0_s1_write;                           // mm_interconnect_0:ram_0_s1_write -> ram_0:write
	wire  [31:0] mm_interconnect_0_ram_0_s1_writedata;                       // mm_interconnect_0:ram_0_s1_writedata -> ram_0:writedata
	wire         mm_interconnect_0_ram_0_s1_clken;                           // mm_interconnect_0:ram_0_s1_clken -> ram_0:clken
	wire  [31:0] mm_interconnect_0_pio_continue_0_s1_readdata;               // pio_continue_0:readdata -> mm_interconnect_0:pio_continue_0_s1_readdata
	wire   [1:0] mm_interconnect_0_pio_continue_0_s1_address;                // mm_interconnect_0:pio_continue_0_s1_address -> pio_continue_0:address
	wire         mm_interconnect_0_pio_leds_0_s1_chipselect;                 // mm_interconnect_0:pio_leds_0_s1_chipselect -> pio_leds_0:chipselect
	wire  [31:0] mm_interconnect_0_pio_leds_0_s1_readdata;                   // pio_leds_0:readdata -> mm_interconnect_0:pio_leds_0_s1_readdata
	wire   [1:0] mm_interconnect_0_pio_leds_0_s1_address;                    // mm_interconnect_0:pio_leds_0_s1_address -> pio_leds_0:address
	wire         mm_interconnect_0_pio_leds_0_s1_write;                      // mm_interconnect_0:pio_leds_0_s1_write -> pio_leds_0:write_n
	wire  [31:0] mm_interconnect_0_pio_leds_0_s1_writedata;                  // mm_interconnect_0:pio_leds_0_s1_writedata -> pio_leds_0:writedata
	wire         mm_interconnect_0_new_sdram_controller_0_s1_chipselect;     // mm_interconnect_0:new_sdram_controller_0_s1_chipselect -> new_sdram_controller_0:az_cs
	wire  [31:0] mm_interconnect_0_new_sdram_controller_0_s1_readdata;       // new_sdram_controller_0:za_data -> mm_interconnect_0:new_sdram_controller_0_s1_readdata
	wire         mm_interconnect_0_new_sdram_controller_0_s1_waitrequest;    // new_sdram_controller_0:za_waitrequest -> mm_interconnect_0:new_sdram_controller_0_s1_waitrequest
	wire  [23:0] mm_interconnect_0_new_sdram_controller_0_s1_address;        // mm_interconnect_0:new_sdram_controller_0_s1_address -> new_sdram_controller_0:az_addr
	wire         mm_interconnect_0_new_sdram_controller_0_s1_read;           // mm_interconnect_0:new_sdram_controller_0_s1_read -> new_sdram_controller_0:az_rd_n
	wire   [3:0] mm_interconnect_0_new_sdram_controller_0_s1_byteenable;     // mm_interconnect_0:new_sdram_controller_0_s1_byteenable -> new_sdram_controller_0:az_be_n
	wire         mm_interconnect_0_new_sdram_controller_0_s1_readdatavalid;  // new_sdram_controller_0:za_valid -> mm_interconnect_0:new_sdram_controller_0_s1_readdatavalid
	wire         mm_interconnect_0_new_sdram_controller_0_s1_write;          // mm_interconnect_0:new_sdram_controller_0_s1_write -> new_sdram_controller_0:az_wr_n
	wire  [31:0] mm_interconnect_0_new_sdram_controller_0_s1_writedata;      // mm_interconnect_0:new_sdram_controller_0_s1_writedata -> new_sdram_controller_0:az_data
	wire         mm_interconnect_0_pio_display1_0_s1_chipselect;             // mm_interconnect_0:pio_display1_0_s1_chipselect -> pio_display1_0:chipselect
	wire  [31:0] mm_interconnect_0_pio_display1_0_s1_readdata;               // pio_display1_0:readdata -> mm_interconnect_0:pio_display1_0_s1_readdata
	wire   [1:0] mm_interconnect_0_pio_display1_0_s1_address;                // mm_interconnect_0:pio_display1_0_s1_address -> pio_display1_0:address
	wire         mm_interconnect_0_pio_display1_0_s1_write;                  // mm_interconnect_0:pio_display1_0_s1_write -> pio_display1_0:write_n
	wire  [31:0] mm_interconnect_0_pio_display1_0_s1_writedata;              // mm_interconnect_0:pio_display1_0_s1_writedata -> pio_display1_0:writedata
	wire         mm_interconnect_0_pio_display2_0_s1_chipselect;             // mm_interconnect_0:pio_display2_0_s1_chipselect -> pio_display2_0:chipselect
	wire  [31:0] mm_interconnect_0_pio_display2_0_s1_readdata;               // pio_display2_0:readdata -> mm_interconnect_0:pio_display2_0_s1_readdata
	wire   [1:0] mm_interconnect_0_pio_display2_0_s1_address;                // mm_interconnect_0:pio_display2_0_s1_address -> pio_display2_0:address
	wire         mm_interconnect_0_pio_display2_0_s1_write;                  // mm_interconnect_0:pio_display2_0_s1_write -> pio_display2_0:write_n
	wire  [31:0] mm_interconnect_0_pio_display2_0_s1_writedata;              // mm_interconnect_0:pio_display2_0_s1_writedata -> pio_display2_0:writedata
	wire         mm_interconnect_0_pio_display3_0_s1_chipselect;             // mm_interconnect_0:pio_display3_0_s1_chipselect -> pio_display3_0:chipselect
	wire  [31:0] mm_interconnect_0_pio_display3_0_s1_readdata;               // pio_display3_0:readdata -> mm_interconnect_0:pio_display3_0_s1_readdata
	wire   [1:0] mm_interconnect_0_pio_display3_0_s1_address;                // mm_interconnect_0:pio_display3_0_s1_address -> pio_display3_0:address
	wire         mm_interconnect_0_pio_display3_0_s1_write;                  // mm_interconnect_0:pio_display3_0_s1_write -> pio_display3_0:write_n
	wire  [31:0] mm_interconnect_0_pio_display3_0_s1_writedata;              // mm_interconnect_0:pio_display3_0_s1_writedata -> pio_display3_0:writedata
	wire         mm_interconnect_0_pio_display4_0_s1_chipselect;             // mm_interconnect_0:pio_display4_0_s1_chipselect -> pio_display4_0:chipselect
	wire  [31:0] mm_interconnect_0_pio_display4_0_s1_readdata;               // pio_display4_0:readdata -> mm_interconnect_0:pio_display4_0_s1_readdata
	wire   [1:0] mm_interconnect_0_pio_display4_0_s1_address;                // mm_interconnect_0:pio_display4_0_s1_address -> pio_display4_0:address
	wire         mm_interconnect_0_pio_display4_0_s1_write;                  // mm_interconnect_0:pio_display4_0_s1_write -> pio_display4_0:write_n
	wire  [31:0] mm_interconnect_0_pio_display4_0_s1_writedata;              // mm_interconnect_0:pio_display4_0_s1_writedata -> pio_display4_0:writedata
	wire         mm_interconnect_0_pio_display5_0_s1_chipselect;             // mm_interconnect_0:pio_display5_0_s1_chipselect -> pio_display5_0:chipselect
	wire  [31:0] mm_interconnect_0_pio_display5_0_s1_readdata;               // pio_display5_0:readdata -> mm_interconnect_0:pio_display5_0_s1_readdata
	wire   [1:0] mm_interconnect_0_pio_display5_0_s1_address;                // mm_interconnect_0:pio_display5_0_s1_address -> pio_display5_0:address
	wire         mm_interconnect_0_pio_display5_0_s1_write;                  // mm_interconnect_0:pio_display5_0_s1_write -> pio_display5_0:write_n
	wire  [31:0] mm_interconnect_0_pio_display5_0_s1_writedata;              // mm_interconnect_0:pio_display5_0_s1_writedata -> pio_display5_0:writedata
	wire         mm_interconnect_0_pio_display6_0_s1_chipselect;             // mm_interconnect_0:pio_display6_0_s1_chipselect -> pio_display6_0:chipselect
	wire  [31:0] mm_interconnect_0_pio_display6_0_s1_readdata;               // pio_display6_0:readdata -> mm_interconnect_0:pio_display6_0_s1_readdata
	wire   [1:0] mm_interconnect_0_pio_display6_0_s1_address;                // mm_interconnect_0:pio_display6_0_s1_address -> pio_display6_0:address
	wire         mm_interconnect_0_pio_display6_0_s1_write;                  // mm_interconnect_0:pio_display6_0_s1_write -> pio_display6_0:write_n
	wire  [31:0] mm_interconnect_0_pio_display6_0_s1_writedata;              // mm_interconnect_0:pio_display6_0_s1_writedata -> pio_display6_0:writedata
	wire  [31:0] mm_interconnect_0_pio_left_right_0_s1_readdata;             // pio_left_right_0:readdata -> mm_interconnect_0:pio_left_right_0_s1_readdata
	wire   [1:0] mm_interconnect_0_pio_left_right_0_s1_address;              // mm_interconnect_0:pio_left_right_0_s1_address -> pio_left_right_0:address
	wire  [31:0] mm_interconnect_0_pio_up_down_0_s1_readdata;                // pio_up_down_0:readdata -> mm_interconnect_0:pio_up_down_0_s1_readdata
	wire   [1:0] mm_interconnect_0_pio_up_down_0_s1_address;                 // mm_interconnect_0:pio_up_down_0_s1_address -> pio_up_down_0:address
	wire         mm_interconnect_0_rom_0_s1_chipselect;                      // mm_interconnect_0:rom_0_s1_chipselect -> rom_0:chipselect
	wire  [31:0] mm_interconnect_0_rom_0_s1_readdata;                        // rom_0:readdata -> mm_interconnect_0:rom_0_s1_readdata
	wire         mm_interconnect_0_rom_0_s1_debugaccess;                     // mm_interconnect_0:rom_0_s1_debugaccess -> rom_0:debugaccess
	wire  [10:0] mm_interconnect_0_rom_0_s1_address;                         // mm_interconnect_0:rom_0_s1_address -> rom_0:address
	wire   [3:0] mm_interconnect_0_rom_0_s1_byteenable;                      // mm_interconnect_0:rom_0_s1_byteenable -> rom_0:byteenable
	wire         mm_interconnect_0_rom_0_s1_write;                           // mm_interconnect_0:rom_0_s1_write -> rom_0:write
	wire  [31:0] mm_interconnect_0_rom_0_s1_writedata;                       // mm_interconnect_0:rom_0_s1_writedata -> rom_0:writedata
	wire         mm_interconnect_0_rom_0_s1_clken;                           // mm_interconnect_0:rom_0_s1_clken -> rom_0:clken
	wire         irq_mapper_receiver0_irq;                                   // timer_0:irq -> irq_mapper:receiver0_irq
	wire  [31:0] nios2_gen2_0_irq_irq;                                       // irq_mapper:sender_irq -> nios2_gen2_0:irq
	wire         rst_controller_reset_out_reset;                             // rst_controller:reset_out -> [irq_mapper:reset, mm_interconnect_0:nios2_gen2_0_reset_reset_bridge_in_reset_reset, new_sdram_controller_0:reset_n, nios2_gen2_0:reset_n, pio_continue_0:reset_n, pio_display1_0:reset_n, pio_display2_0:reset_n, pio_display3_0:reset_n, pio_display4_0:reset_n, pio_display5_0:reset_n, pio_display6_0:reset_n, pio_leds_0:reset_n, pio_left_right_0:reset_n, pio_up_down_0:reset_n, ram_0:reset, rom_0:reset, rst_translator:in_reset, timer_0:reset_n]
	wire         rst_controller_reset_out_reset_req;                         // rst_controller:reset_req -> [nios2_gen2_0:reset_req, ram_0:reset_req, rom_0:reset_req, rst_translator:reset_req_in]

	cpuqsys_new_sdram_controller_0 new_sdram_controller_0 (
		.clk            (clk_clk),                                                   //   clk.clk
		.reset_n        (~rst_controller_reset_out_reset),                           // reset.reset_n
		.az_addr        (mm_interconnect_0_new_sdram_controller_0_s1_address),       //    s1.address
		.az_be_n        (~mm_interconnect_0_new_sdram_controller_0_s1_byteenable),   //      .byteenable_n
		.az_cs          (mm_interconnect_0_new_sdram_controller_0_s1_chipselect),    //      .chipselect
		.az_data        (mm_interconnect_0_new_sdram_controller_0_s1_writedata),     //      .writedata
		.az_rd_n        (~mm_interconnect_0_new_sdram_controller_0_s1_read),         //      .read_n
		.az_wr_n        (~mm_interconnect_0_new_sdram_controller_0_s1_write),        //      .write_n
		.za_data        (mm_interconnect_0_new_sdram_controller_0_s1_readdata),      //      .readdata
		.za_valid       (mm_interconnect_0_new_sdram_controller_0_s1_readdatavalid), //      .readdatavalid
		.za_waitrequest (mm_interconnect_0_new_sdram_controller_0_s1_waitrequest),   //      .waitrequest
		.zs_addr        (new_sdram_controller_0_wire_addr),                          //  wire.export
		.zs_ba          (new_sdram_controller_0_wire_ba),                            //      .export
		.zs_cas_n       (new_sdram_controller_0_wire_cas_n),                         //      .export
		.zs_cke         (new_sdram_controller_0_wire_cke),                           //      .export
		.zs_cs_n        (new_sdram_controller_0_wire_cs_n),                          //      .export
		.zs_dq          (new_sdram_controller_0_wire_dq),                            //      .export
		.zs_dqm         (new_sdram_controller_0_wire_dqm),                           //      .export
		.zs_ras_n       (new_sdram_controller_0_wire_ras_n),                         //      .export
		.zs_we_n        (new_sdram_controller_0_wire_we_n)                           //      .export
	);

	cpuqsys_nios2_gen2_0 nios2_gen2_0 (
		.clk                                 (clk_clk),                                                    //                       clk.clk
		.reset_n                             (~rst_controller_reset_out_reset),                            //                     reset.reset_n
		.reset_req                           (rst_controller_reset_out_reset_req),                         //                          .reset_req
		.d_address                           (nios2_gen2_0_data_master_address),                           //               data_master.address
		.d_byteenable                        (nios2_gen2_0_data_master_byteenable),                        //                          .byteenable
		.d_read                              (nios2_gen2_0_data_master_read),                              //                          .read
		.d_readdata                          (nios2_gen2_0_data_master_readdata),                          //                          .readdata
		.d_waitrequest                       (nios2_gen2_0_data_master_waitrequest),                       //                          .waitrequest
		.d_write                             (nios2_gen2_0_data_master_write),                             //                          .write
		.d_writedata                         (nios2_gen2_0_data_master_writedata),                         //                          .writedata
		.debug_mem_slave_debugaccess_to_roms (nios2_gen2_0_data_master_debugaccess),                       //                          .debugaccess
		.i_address                           (nios2_gen2_0_instruction_master_address),                    //        instruction_master.address
		.i_read                              (nios2_gen2_0_instruction_master_read),                       //                          .read
		.i_readdata                          (nios2_gen2_0_instruction_master_readdata),                   //                          .readdata
		.i_waitrequest                       (nios2_gen2_0_instruction_master_waitrequest),                //                          .waitrequest
		.irq                                 (nios2_gen2_0_irq_irq),                                       //                       irq.irq
		.debug_reset_request                 (),                                                           //       debug_reset_request.reset
		.debug_mem_slave_address             (mm_interconnect_0_nios2_gen2_0_debug_mem_slave_address),     //           debug_mem_slave.address
		.debug_mem_slave_byteenable          (mm_interconnect_0_nios2_gen2_0_debug_mem_slave_byteenable),  //                          .byteenable
		.debug_mem_slave_debugaccess         (mm_interconnect_0_nios2_gen2_0_debug_mem_slave_debugaccess), //                          .debugaccess
		.debug_mem_slave_read                (mm_interconnect_0_nios2_gen2_0_debug_mem_slave_read),        //                          .read
		.debug_mem_slave_readdata            (mm_interconnect_0_nios2_gen2_0_debug_mem_slave_readdata),    //                          .readdata
		.debug_mem_slave_waitrequest         (mm_interconnect_0_nios2_gen2_0_debug_mem_slave_waitrequest), //                          .waitrequest
		.debug_mem_slave_write               (mm_interconnect_0_nios2_gen2_0_debug_mem_slave_write),       //                          .write
		.debug_mem_slave_writedata           (mm_interconnect_0_nios2_gen2_0_debug_mem_slave_writedata),   //                          .writedata
		.dummy_ci_port                       ()                                                            // custom_instruction_master.readra
	);

	cpuqsys_pio_continue_0 pio_continue_0 (
		.clk      (clk_clk),                                      //                 clk.clk
		.reset_n  (~rst_controller_reset_out_reset),              //               reset.reset_n
		.address  (mm_interconnect_0_pio_continue_0_s1_address),  //                  s1.address
		.readdata (mm_interconnect_0_pio_continue_0_s1_readdata), //                    .readdata
		.in_port  (pio_continue_0_external_connection_export)     // external_connection.export
	);

	cpuqsys_pio_display1_0 pio_display1_0 (
		.clk        (clk_clk),                                        //                 clk.clk
		.reset_n    (~rst_controller_reset_out_reset),                //               reset.reset_n
		.address    (mm_interconnect_0_pio_display1_0_s1_address),    //                  s1.address
		.write_n    (~mm_interconnect_0_pio_display1_0_s1_write),     //                    .write_n
		.writedata  (mm_interconnect_0_pio_display1_0_s1_writedata),  //                    .writedata
		.chipselect (mm_interconnect_0_pio_display1_0_s1_chipselect), //                    .chipselect
		.readdata   (mm_interconnect_0_pio_display1_0_s1_readdata),   //                    .readdata
		.out_port   (pio_display1_0_external_connection_export)       // external_connection.export
	);

	cpuqsys_pio_display1_0 pio_display2_0 (
		.clk        (clk_clk),                                        //                 clk.clk
		.reset_n    (~rst_controller_reset_out_reset),                //               reset.reset_n
		.address    (mm_interconnect_0_pio_display2_0_s1_address),    //                  s1.address
		.write_n    (~mm_interconnect_0_pio_display2_0_s1_write),     //                    .write_n
		.writedata  (mm_interconnect_0_pio_display2_0_s1_writedata),  //                    .writedata
		.chipselect (mm_interconnect_0_pio_display2_0_s1_chipselect), //                    .chipselect
		.readdata   (mm_interconnect_0_pio_display2_0_s1_readdata),   //                    .readdata
		.out_port   (pio_display2_0_external_connection_export)       // external_connection.export
	);

	cpuqsys_pio_display1_0 pio_display3_0 (
		.clk        (clk_clk),                                        //                 clk.clk
		.reset_n    (~rst_controller_reset_out_reset),                //               reset.reset_n
		.address    (mm_interconnect_0_pio_display3_0_s1_address),    //                  s1.address
		.write_n    (~mm_interconnect_0_pio_display3_0_s1_write),     //                    .write_n
		.writedata  (mm_interconnect_0_pio_display3_0_s1_writedata),  //                    .writedata
		.chipselect (mm_interconnect_0_pio_display3_0_s1_chipselect), //                    .chipselect
		.readdata   (mm_interconnect_0_pio_display3_0_s1_readdata),   //                    .readdata
		.out_port   (pio_display3_0_external_connection_export)       // external_connection.export
	);

	cpuqsys_pio_display1_0 pio_display4_0 (
		.clk        (clk_clk),                                        //                 clk.clk
		.reset_n    (~rst_controller_reset_out_reset),                //               reset.reset_n
		.address    (mm_interconnect_0_pio_display4_0_s1_address),    //                  s1.address
		.write_n    (~mm_interconnect_0_pio_display4_0_s1_write),     //                    .write_n
		.writedata  (mm_interconnect_0_pio_display4_0_s1_writedata),  //                    .writedata
		.chipselect (mm_interconnect_0_pio_display4_0_s1_chipselect), //                    .chipselect
		.readdata   (mm_interconnect_0_pio_display4_0_s1_readdata),   //                    .readdata
		.out_port   (pio_display4_0_external_connection_export)       // external_connection.export
	);

	cpuqsys_pio_display1_0 pio_display5_0 (
		.clk        (clk_clk),                                        //                 clk.clk
		.reset_n    (~rst_controller_reset_out_reset),                //               reset.reset_n
		.address    (mm_interconnect_0_pio_display5_0_s1_address),    //                  s1.address
		.write_n    (~mm_interconnect_0_pio_display5_0_s1_write),     //                    .write_n
		.writedata  (mm_interconnect_0_pio_display5_0_s1_writedata),  //                    .writedata
		.chipselect (mm_interconnect_0_pio_display5_0_s1_chipselect), //                    .chipselect
		.readdata   (mm_interconnect_0_pio_display5_0_s1_readdata),   //                    .readdata
		.out_port   (pio_display5_0_external_connection_export)       // external_connection.export
	);

	cpuqsys_pio_display1_0 pio_display6_0 (
		.clk        (clk_clk),                                        //                 clk.clk
		.reset_n    (~rst_controller_reset_out_reset),                //               reset.reset_n
		.address    (mm_interconnect_0_pio_display6_0_s1_address),    //                  s1.address
		.write_n    (~mm_interconnect_0_pio_display6_0_s1_write),     //                    .write_n
		.writedata  (mm_interconnect_0_pio_display6_0_s1_writedata),  //                    .writedata
		.chipselect (mm_interconnect_0_pio_display6_0_s1_chipselect), //                    .chipselect
		.readdata   (mm_interconnect_0_pio_display6_0_s1_readdata),   //                    .readdata
		.out_port   (pio_display6_0_external_connection_export)       // external_connection.export
	);

	cpuqsys_pio_leds_0 pio_leds_0 (
		.clk        (clk_clk),                                    //                 clk.clk
		.reset_n    (~rst_controller_reset_out_reset),            //               reset.reset_n
		.address    (mm_interconnect_0_pio_leds_0_s1_address),    //                  s1.address
		.write_n    (~mm_interconnect_0_pio_leds_0_s1_write),     //                    .write_n
		.writedata  (mm_interconnect_0_pio_leds_0_s1_writedata),  //                    .writedata
		.chipselect (mm_interconnect_0_pio_leds_0_s1_chipselect), //                    .chipselect
		.readdata   (mm_interconnect_0_pio_leds_0_s1_readdata),   //                    .readdata
		.out_port   (pio_leds_0_external_connection_export)       // external_connection.export
	);

	cpuqsys_pio_left_right_0 pio_left_right_0 (
		.clk      (clk_clk),                                        //                 clk.clk
		.reset_n  (~rst_controller_reset_out_reset),                //               reset.reset_n
		.address  (mm_interconnect_0_pio_left_right_0_s1_address),  //                  s1.address
		.readdata (mm_interconnect_0_pio_left_right_0_s1_readdata), //                    .readdata
		.in_port  (pio_left_right_0_external_connection_export)     // external_connection.export
	);

	cpuqsys_pio_left_right_0 pio_up_down_0 (
		.clk      (clk_clk),                                     //                 clk.clk
		.reset_n  (~rst_controller_reset_out_reset),             //               reset.reset_n
		.address  (mm_interconnect_0_pio_up_down_0_s1_address),  //                  s1.address
		.readdata (mm_interconnect_0_pio_up_down_0_s1_readdata), //                    .readdata
		.in_port  (pio_up_down_0_external_connection_export)     // external_connection.export
	);

	cpuqsys_ram_0 ram_0 (
		.clk        (clk_clk),                               //   clk1.clk
		.address    (mm_interconnect_0_ram_0_s1_address),    //     s1.address
		.clken      (mm_interconnect_0_ram_0_s1_clken),      //       .clken
		.chipselect (mm_interconnect_0_ram_0_s1_chipselect), //       .chipselect
		.write      (mm_interconnect_0_ram_0_s1_write),      //       .write
		.readdata   (mm_interconnect_0_ram_0_s1_readdata),   //       .readdata
		.writedata  (mm_interconnect_0_ram_0_s1_writedata),  //       .writedata
		.byteenable (mm_interconnect_0_ram_0_s1_byteenable), //       .byteenable
		.reset      (rst_controller_reset_out_reset),        // reset1.reset
		.reset_req  (rst_controller_reset_out_reset_req),    //       .reset_req
		.freeze     (1'b0)                                   // (terminated)
	);

	cpuqsys_rom_0 rom_0 (
		.clk         (clk_clk),                                //   clk1.clk
		.address     (mm_interconnect_0_rom_0_s1_address),     //     s1.address
		.debugaccess (mm_interconnect_0_rom_0_s1_debugaccess), //       .debugaccess
		.clken       (mm_interconnect_0_rom_0_s1_clken),       //       .clken
		.chipselect  (mm_interconnect_0_rom_0_s1_chipselect),  //       .chipselect
		.write       (mm_interconnect_0_rom_0_s1_write),       //       .write
		.readdata    (mm_interconnect_0_rom_0_s1_readdata),    //       .readdata
		.writedata   (mm_interconnect_0_rom_0_s1_writedata),   //       .writedata
		.byteenable  (mm_interconnect_0_rom_0_s1_byteenable),  //       .byteenable
		.reset       (rst_controller_reset_out_reset),         // reset1.reset
		.reset_req   (rst_controller_reset_out_reset_req),     //       .reset_req
		.freeze      (1'b0)                                    // (terminated)
	);

	cpuqsys_timer_0 timer_0 (
		.clk        (clk_clk),                                 //   clk.clk
		.reset_n    (~rst_controller_reset_out_reset),         // reset.reset_n
		.address    (mm_interconnect_0_timer_0_s1_address),    //    s1.address
		.writedata  (mm_interconnect_0_timer_0_s1_writedata),  //      .writedata
		.readdata   (mm_interconnect_0_timer_0_s1_readdata),   //      .readdata
		.chipselect (mm_interconnect_0_timer_0_s1_chipselect), //      .chipselect
		.write_n    (~mm_interconnect_0_timer_0_s1_write),     //      .write_n
		.irq        (irq_mapper_receiver0_irq)                 //   irq.irq
	);

	cpuqsys_mm_interconnect_0 mm_interconnect_0 (
		.clk_0_clk_clk                                  (clk_clk),                                                    //                                clk_0_clk.clk
		.nios2_gen2_0_reset_reset_bridge_in_reset_reset (rst_controller_reset_out_reset),                             // nios2_gen2_0_reset_reset_bridge_in_reset.reset
		.nios2_gen2_0_data_master_address               (nios2_gen2_0_data_master_address),                           //                 nios2_gen2_0_data_master.address
		.nios2_gen2_0_data_master_waitrequest           (nios2_gen2_0_data_master_waitrequest),                       //                                         .waitrequest
		.nios2_gen2_0_data_master_byteenable            (nios2_gen2_0_data_master_byteenable),                        //                                         .byteenable
		.nios2_gen2_0_data_master_read                  (nios2_gen2_0_data_master_read),                              //                                         .read
		.nios2_gen2_0_data_master_readdata              (nios2_gen2_0_data_master_readdata),                          //                                         .readdata
		.nios2_gen2_0_data_master_write                 (nios2_gen2_0_data_master_write),                             //                                         .write
		.nios2_gen2_0_data_master_writedata             (nios2_gen2_0_data_master_writedata),                         //                                         .writedata
		.nios2_gen2_0_data_master_debugaccess           (nios2_gen2_0_data_master_debugaccess),                       //                                         .debugaccess
		.nios2_gen2_0_instruction_master_address        (nios2_gen2_0_instruction_master_address),                    //          nios2_gen2_0_instruction_master.address
		.nios2_gen2_0_instruction_master_waitrequest    (nios2_gen2_0_instruction_master_waitrequest),                //                                         .waitrequest
		.nios2_gen2_0_instruction_master_read           (nios2_gen2_0_instruction_master_read),                       //                                         .read
		.nios2_gen2_0_instruction_master_readdata       (nios2_gen2_0_instruction_master_readdata),                   //                                         .readdata
		.new_sdram_controller_0_s1_address              (mm_interconnect_0_new_sdram_controller_0_s1_address),        //                new_sdram_controller_0_s1.address
		.new_sdram_controller_0_s1_write                (mm_interconnect_0_new_sdram_controller_0_s1_write),          //                                         .write
		.new_sdram_controller_0_s1_read                 (mm_interconnect_0_new_sdram_controller_0_s1_read),           //                                         .read
		.new_sdram_controller_0_s1_readdata             (mm_interconnect_0_new_sdram_controller_0_s1_readdata),       //                                         .readdata
		.new_sdram_controller_0_s1_writedata            (mm_interconnect_0_new_sdram_controller_0_s1_writedata),      //                                         .writedata
		.new_sdram_controller_0_s1_byteenable           (mm_interconnect_0_new_sdram_controller_0_s1_byteenable),     //                                         .byteenable
		.new_sdram_controller_0_s1_readdatavalid        (mm_interconnect_0_new_sdram_controller_0_s1_readdatavalid),  //                                         .readdatavalid
		.new_sdram_controller_0_s1_waitrequest          (mm_interconnect_0_new_sdram_controller_0_s1_waitrequest),    //                                         .waitrequest
		.new_sdram_controller_0_s1_chipselect           (mm_interconnect_0_new_sdram_controller_0_s1_chipselect),     //                                         .chipselect
		.nios2_gen2_0_debug_mem_slave_address           (mm_interconnect_0_nios2_gen2_0_debug_mem_slave_address),     //             nios2_gen2_0_debug_mem_slave.address
		.nios2_gen2_0_debug_mem_slave_write             (mm_interconnect_0_nios2_gen2_0_debug_mem_slave_write),       //                                         .write
		.nios2_gen2_0_debug_mem_slave_read              (mm_interconnect_0_nios2_gen2_0_debug_mem_slave_read),        //                                         .read
		.nios2_gen2_0_debug_mem_slave_readdata          (mm_interconnect_0_nios2_gen2_0_debug_mem_slave_readdata),    //                                         .readdata
		.nios2_gen2_0_debug_mem_slave_writedata         (mm_interconnect_0_nios2_gen2_0_debug_mem_slave_writedata),   //                                         .writedata
		.nios2_gen2_0_debug_mem_slave_byteenable        (mm_interconnect_0_nios2_gen2_0_debug_mem_slave_byteenable),  //                                         .byteenable
		.nios2_gen2_0_debug_mem_slave_waitrequest       (mm_interconnect_0_nios2_gen2_0_debug_mem_slave_waitrequest), //                                         .waitrequest
		.nios2_gen2_0_debug_mem_slave_debugaccess       (mm_interconnect_0_nios2_gen2_0_debug_mem_slave_debugaccess), //                                         .debugaccess
		.pio_continue_0_s1_address                      (mm_interconnect_0_pio_continue_0_s1_address),                //                        pio_continue_0_s1.address
		.pio_continue_0_s1_readdata                     (mm_interconnect_0_pio_continue_0_s1_readdata),               //                                         .readdata
		.pio_display1_0_s1_address                      (mm_interconnect_0_pio_display1_0_s1_address),                //                        pio_display1_0_s1.address
		.pio_display1_0_s1_write                        (mm_interconnect_0_pio_display1_0_s1_write),                  //                                         .write
		.pio_display1_0_s1_readdata                     (mm_interconnect_0_pio_display1_0_s1_readdata),               //                                         .readdata
		.pio_display1_0_s1_writedata                    (mm_interconnect_0_pio_display1_0_s1_writedata),              //                                         .writedata
		.pio_display1_0_s1_chipselect                   (mm_interconnect_0_pio_display1_0_s1_chipselect),             //                                         .chipselect
		.pio_display2_0_s1_address                      (mm_interconnect_0_pio_display2_0_s1_address),                //                        pio_display2_0_s1.address
		.pio_display2_0_s1_write                        (mm_interconnect_0_pio_display2_0_s1_write),                  //                                         .write
		.pio_display2_0_s1_readdata                     (mm_interconnect_0_pio_display2_0_s1_readdata),               //                                         .readdata
		.pio_display2_0_s1_writedata                    (mm_interconnect_0_pio_display2_0_s1_writedata),              //                                         .writedata
		.pio_display2_0_s1_chipselect                   (mm_interconnect_0_pio_display2_0_s1_chipselect),             //                                         .chipselect
		.pio_display3_0_s1_address                      (mm_interconnect_0_pio_display3_0_s1_address),                //                        pio_display3_0_s1.address
		.pio_display3_0_s1_write                        (mm_interconnect_0_pio_display3_0_s1_write),                  //                                         .write
		.pio_display3_0_s1_readdata                     (mm_interconnect_0_pio_display3_0_s1_readdata),               //                                         .readdata
		.pio_display3_0_s1_writedata                    (mm_interconnect_0_pio_display3_0_s1_writedata),              //                                         .writedata
		.pio_display3_0_s1_chipselect                   (mm_interconnect_0_pio_display3_0_s1_chipselect),             //                                         .chipselect
		.pio_display4_0_s1_address                      (mm_interconnect_0_pio_display4_0_s1_address),                //                        pio_display4_0_s1.address
		.pio_display4_0_s1_write                        (mm_interconnect_0_pio_display4_0_s1_write),                  //                                         .write
		.pio_display4_0_s1_readdata                     (mm_interconnect_0_pio_display4_0_s1_readdata),               //                                         .readdata
		.pio_display4_0_s1_writedata                    (mm_interconnect_0_pio_display4_0_s1_writedata),              //                                         .writedata
		.pio_display4_0_s1_chipselect                   (mm_interconnect_0_pio_display4_0_s1_chipselect),             //                                         .chipselect
		.pio_display5_0_s1_address                      (mm_interconnect_0_pio_display5_0_s1_address),                //                        pio_display5_0_s1.address
		.pio_display5_0_s1_write                        (mm_interconnect_0_pio_display5_0_s1_write),                  //                                         .write
		.pio_display5_0_s1_readdata                     (mm_interconnect_0_pio_display5_0_s1_readdata),               //                                         .readdata
		.pio_display5_0_s1_writedata                    (mm_interconnect_0_pio_display5_0_s1_writedata),              //                                         .writedata
		.pio_display5_0_s1_chipselect                   (mm_interconnect_0_pio_display5_0_s1_chipselect),             //                                         .chipselect
		.pio_display6_0_s1_address                      (mm_interconnect_0_pio_display6_0_s1_address),                //                        pio_display6_0_s1.address
		.pio_display6_0_s1_write                        (mm_interconnect_0_pio_display6_0_s1_write),                  //                                         .write
		.pio_display6_0_s1_readdata                     (mm_interconnect_0_pio_display6_0_s1_readdata),               //                                         .readdata
		.pio_display6_0_s1_writedata                    (mm_interconnect_0_pio_display6_0_s1_writedata),              //                                         .writedata
		.pio_display6_0_s1_chipselect                   (mm_interconnect_0_pio_display6_0_s1_chipselect),             //                                         .chipselect
		.pio_leds_0_s1_address                          (mm_interconnect_0_pio_leds_0_s1_address),                    //                            pio_leds_0_s1.address
		.pio_leds_0_s1_write                            (mm_interconnect_0_pio_leds_0_s1_write),                      //                                         .write
		.pio_leds_0_s1_readdata                         (mm_interconnect_0_pio_leds_0_s1_readdata),                   //                                         .readdata
		.pio_leds_0_s1_writedata                        (mm_interconnect_0_pio_leds_0_s1_writedata),                  //                                         .writedata
		.pio_leds_0_s1_chipselect                       (mm_interconnect_0_pio_leds_0_s1_chipselect),                 //                                         .chipselect
		.pio_left_right_0_s1_address                    (mm_interconnect_0_pio_left_right_0_s1_address),              //                      pio_left_right_0_s1.address
		.pio_left_right_0_s1_readdata                   (mm_interconnect_0_pio_left_right_0_s1_readdata),             //                                         .readdata
		.pio_up_down_0_s1_address                       (mm_interconnect_0_pio_up_down_0_s1_address),                 //                         pio_up_down_0_s1.address
		.pio_up_down_0_s1_readdata                      (mm_interconnect_0_pio_up_down_0_s1_readdata),                //                                         .readdata
		.ram_0_s1_address                               (mm_interconnect_0_ram_0_s1_address),                         //                                 ram_0_s1.address
		.ram_0_s1_write                                 (mm_interconnect_0_ram_0_s1_write),                           //                                         .write
		.ram_0_s1_readdata                              (mm_interconnect_0_ram_0_s1_readdata),                        //                                         .readdata
		.ram_0_s1_writedata                             (mm_interconnect_0_ram_0_s1_writedata),                       //                                         .writedata
		.ram_0_s1_byteenable                            (mm_interconnect_0_ram_0_s1_byteenable),                      //                                         .byteenable
		.ram_0_s1_chipselect                            (mm_interconnect_0_ram_0_s1_chipselect),                      //                                         .chipselect
		.ram_0_s1_clken                                 (mm_interconnect_0_ram_0_s1_clken),                           //                                         .clken
		.rom_0_s1_address                               (mm_interconnect_0_rom_0_s1_address),                         //                                 rom_0_s1.address
		.rom_0_s1_write                                 (mm_interconnect_0_rom_0_s1_write),                           //                                         .write
		.rom_0_s1_readdata                              (mm_interconnect_0_rom_0_s1_readdata),                        //                                         .readdata
		.rom_0_s1_writedata                             (mm_interconnect_0_rom_0_s1_writedata),                       //                                         .writedata
		.rom_0_s1_byteenable                            (mm_interconnect_0_rom_0_s1_byteenable),                      //                                         .byteenable
		.rom_0_s1_chipselect                            (mm_interconnect_0_rom_0_s1_chipselect),                      //                                         .chipselect
		.rom_0_s1_clken                                 (mm_interconnect_0_rom_0_s1_clken),                           //                                         .clken
		.rom_0_s1_debugaccess                           (mm_interconnect_0_rom_0_s1_debugaccess),                     //                                         .debugaccess
		.timer_0_s1_address                             (mm_interconnect_0_timer_0_s1_address),                       //                               timer_0_s1.address
		.timer_0_s1_write                               (mm_interconnect_0_timer_0_s1_write),                         //                                         .write
		.timer_0_s1_readdata                            (mm_interconnect_0_timer_0_s1_readdata),                      //                                         .readdata
		.timer_0_s1_writedata                           (mm_interconnect_0_timer_0_s1_writedata),                     //                                         .writedata
		.timer_0_s1_chipselect                          (mm_interconnect_0_timer_0_s1_chipselect)                     //                                         .chipselect
	);

	cpuqsys_irq_mapper irq_mapper (
		.clk           (clk_clk),                        //       clk.clk
		.reset         (rst_controller_reset_out_reset), // clk_reset.reset
		.receiver0_irq (irq_mapper_receiver0_irq),       // receiver0.irq
		.sender_irq    (nios2_gen2_0_irq_irq)            //    sender.irq
	);

	altera_reset_controller #(
		.NUM_RESET_INPUTS          (1),
		.OUTPUT_RESET_SYNC_EDGES   ("deassert"),
		.SYNC_DEPTH                (2),
		.RESET_REQUEST_PRESENT     (1),
		.RESET_REQ_WAIT_TIME       (1),
		.MIN_RST_ASSERTION_TIME    (3),
		.RESET_REQ_EARLY_DSRT_TIME (1),
		.USE_RESET_REQUEST_IN0     (0),
		.USE_RESET_REQUEST_IN1     (0),
		.USE_RESET_REQUEST_IN2     (0),
		.USE_RESET_REQUEST_IN3     (0),
		.USE_RESET_REQUEST_IN4     (0),
		.USE_RESET_REQUEST_IN5     (0),
		.USE_RESET_REQUEST_IN6     (0),
		.USE_RESET_REQUEST_IN7     (0),
		.USE_RESET_REQUEST_IN8     (0),
		.USE_RESET_REQUEST_IN9     (0),
		.USE_RESET_REQUEST_IN10    (0),
		.USE_RESET_REQUEST_IN11    (0),
		.USE_RESET_REQUEST_IN12    (0),
		.USE_RESET_REQUEST_IN13    (0),
		.USE_RESET_REQUEST_IN14    (0),
		.USE_RESET_REQUEST_IN15    (0),
		.ADAPT_RESET_REQUEST       (0)
	) rst_controller (
		.reset_in0      (~reset_reset_n),                     // reset_in0.reset
		.clk            (clk_clk),                            //       clk.clk
		.reset_out      (rst_controller_reset_out_reset),     // reset_out.reset
		.reset_req      (rst_controller_reset_out_reset_req), //          .reset_req
		.reset_req_in0  (1'b0),                               // (terminated)
		.reset_in1      (1'b0),                               // (terminated)
		.reset_req_in1  (1'b0),                               // (terminated)
		.reset_in2      (1'b0),                               // (terminated)
		.reset_req_in2  (1'b0),                               // (terminated)
		.reset_in3      (1'b0),                               // (terminated)
		.reset_req_in3  (1'b0),                               // (terminated)
		.reset_in4      (1'b0),                               // (terminated)
		.reset_req_in4  (1'b0),                               // (terminated)
		.reset_in5      (1'b0),                               // (terminated)
		.reset_req_in5  (1'b0),                               // (terminated)
		.reset_in6      (1'b0),                               // (terminated)
		.reset_req_in6  (1'b0),                               // (terminated)
		.reset_in7      (1'b0),                               // (terminated)
		.reset_req_in7  (1'b0),                               // (terminated)
		.reset_in8      (1'b0),                               // (terminated)
		.reset_req_in8  (1'b0),                               // (terminated)
		.reset_in9      (1'b0),                               // (terminated)
		.reset_req_in9  (1'b0),                               // (terminated)
		.reset_in10     (1'b0),                               // (terminated)
		.reset_req_in10 (1'b0),                               // (terminated)
		.reset_in11     (1'b0),                               // (terminated)
		.reset_req_in11 (1'b0),                               // (terminated)
		.reset_in12     (1'b0),                               // (terminated)
		.reset_req_in12 (1'b0),                               // (terminated)
		.reset_in13     (1'b0),                               // (terminated)
		.reset_req_in13 (1'b0),                               // (terminated)
		.reset_in14     (1'b0),                               // (terminated)
		.reset_req_in14 (1'b0),                               // (terminated)
		.reset_in15     (1'b0),                               // (terminated)
		.reset_req_in15 (1'b0)                                // (terminated)
	);

endmodule
